-- MUX_MEM_WB.vhd

ENTITY MUX_MEM_WB IS 
END MUX_MEM_WB;

ARCHITECTURE Behaviour OF MUX_MEM_WB IS

BEGIN


END Behaviour;