-- MUX_EXE_MEM.vhd

ENTITY MUX_EXE_MEM IS
END MUX_EXE_MEM;

ARCHITECTURE Behaviour OF MUX_EXE_MEM IS

BEGIN


END Behaviour;