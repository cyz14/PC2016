-- DataMemory.vhd

ENTITY DataMemory IS PORT (
    IN     STD_LOGIC;
    IN     STD_LOGIC_VECTOR;
    OUT    STD_LOGIC;
    OUT    STD_LOGIC_VECTOR
);
END DataMemory;

ARCHITECTURE Behaviour OF DataMemory IS

BEGIN


END Behaviour;