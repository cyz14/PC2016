
ENTITY Ctrl_WB IS PORT (

);
END Ctrl_WB;
