-- BubbleStallUnit

ENTITY BubbleStallUnit IS
PORT (
    CLK      :  IN     STD_LOGIC
);
END BubbleStallUnit;


ARCHITECTURE Behaviour OF BubbleStallUnit IS

BEGIN


END Behaviour;