-- MUX_ID_EXE.vhd

ENTITY MUX_ID_EXE IS PORT (
    IN     STD_LOGIC;
    IN     STD_LOGIC_VECTOR;
    OUT    STD_LOGIC;
    OUT    STD_LOGIC_VECTOR
);
END MUX_ID_EXE;

ARCHITECTURE Behaviour OF MUX_ID_EXE IS

BEGIN


END Behaviour;