-- MUX_MEM_WB.vhd

ENTITY MUX_MEM_WB IS PORT (
    IN     STD_LOGIC;
    IN     STD_LOGIC_VECTOR;
    OUT    STD_LOGIC;
    OUT    STD_LOGIC_VECTOR
);
END MUX_MEM_WB;

ARCHITECTURE Behaviour OF MUX_MEM_WB IS

BEGIN


END Behaviour;