ENTITY Ctrl_M IS PORT (
    
);
END Ctrl_M;