-- MUX_EXE_MEM.vhd

ENTITY MUX_EXE_MEM IS PORT (
    IN     STD_LOGIC;
    IN     STD_LOGIC_VECTOR;
    OUT    STD_LOGIC;
    OUT    STD_LOGIC_VECTOR
);
END MUX_EXE_MEM;

ARCHITECTURE Behaviour OF MUX_EXE_MEM IS

BEGIN


END Behaviour;