-- BubbleStallUnit

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY BubbleStallUnit IS
PORT (
    CLK      :  IN     STD_LOGIC
);
END BubbleStallUnit;


ARCHITECTURE Behaviour OF BubbleStallUnit IS

BEGIN


END Behaviour;